library ieee; 
USE ieee.std_logic_1164.all;

entity Save_Register is
end Save_Register;

architecture behaviour of Save_Register